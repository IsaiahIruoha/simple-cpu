module encoder_32_to_5 (input wire [31:0] encoderInput, output reg [4:0] encoderOutput);
	always @ (*) begin
    case (encoderInput)
        32'b00000000000000000000000000000001: encoderOutput <= 5'd0;
		  32'b00000000000000000000000000000010: encoderOutput <= 5'd1;
		  32'b00000000000000000000000000000100: encoderOutput <= 5'd2;
		  32'b00000000000000000000000000001000: encoderOutput <= 5'd3;
		  32'b00000000000000000000000000010000: encoderOutput <= 5'd4;
		  32'b00000000000000000000000000100000: encoderOutput <= 5'd5;
		  32'b00000000000000000000000001000000: encoderOutput <= 5'd6;
		  32'b00000000000000000000000010000000: encoderOutput <= 5'd7;
		  32'b00000000000000000000000100000000: encoderOutput <= 5'd8;
		  32'b00000000000000000000001000000000: encoderOutput <= 5'd9;
		  32'b00000000000000000000010000000000: encoderOutput <= 5'd10;
		  32'b00000000000000000000100000000000: encoderOutput <= 5'd11;
		  32'b00000000000000000001000000000000: encoderOutput <= 5'd12;
		  32'b00000000000000000010000000000000: encoderOutput <= 5'd13;
		  32'b00000000000000000100000000000000: encoderOutput <= 5'd14;
		  32'b00000000000000001000000000000000: encoderOutput <= 5'd15;
		  32'b00000000000000010000000000000000: encoderOutput <= 5'd16;
		  32'b00000000000000100000000000000000: encoderOutput <= 5'd17;
		  32'b00000000000001000000000000000000: encoderOutput <= 5'd18;
		  32'b00000000000010000000000000000000: encoderOutput <= 5'd19;
		  32'b00000000000100000000000000000000: encoderOutput <= 5'd20;
		  32'b00000000001000000000000000000000: encoderOutput <= 5'd21;
		  32'b00000000010000000000000000000000: encoderOutput <= 5'd22;
		  32'b00000000100000000000000000000000: encoderOutput <= 5'd23;   
        default: encoderOutput <= 5'd31;
    endcase
	end
endmodule
